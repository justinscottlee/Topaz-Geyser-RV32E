`timescale 1ns / 1ps

module topaz_geyser_core(
    input logic clk, rst
    );
    
    
    
endmodule